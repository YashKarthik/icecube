`default_nettype none

module main (
    input wire clk
);
endmodule
