`default_nettype none

module matmul (
    input wire i_clk,
    input wire i_trigger,
    input wire i_m,
    input wire i_n
);
endmodule
